module ethernet_test_top ();

endmodule
