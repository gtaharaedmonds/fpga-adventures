module ethernet_test_top ();
  axi_ethernetlite_0 axi_ethernetlite_inst ();
endmodule
